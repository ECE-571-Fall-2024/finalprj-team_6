module M_PC_ADDER(input logic [31:0] a, b, output[31:0] y);
    assign y = a + b;
endmodule